`define CYCLE_TIME 20
`define INSTRUCTION_NUMBERS 500		//此行修改INSTRUCTION_NUMBERS
`timescale 1ns/1ps
`include "CPU.v"

module testbench;
reg Clk, Rst;
reg [31:0] cycles, i;

// Instruction DM initialilation
initial
begin
	/*=================================================     write down your program     =================================================*/


cpu.IF.instruction[0] = 32'b100011_00000_01000_0000000000000000;	//lw r8, r0, 0
cpu.IF.instruction[1] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[2] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[3] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[4] = 32'b000000_00000_00000_10011_00000_100000;	//add r19, r0, r0
cpu.IF.instruction[5] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[6] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[7] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[8] = 32'b000100_01000_00011_00000_00000_000111;	//beq r8, r3, ,special_3
cpu.IF.instruction[9] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[10] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[11] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[12] = 32'b000010_00000_00000_00000_00000_011100;	//j non_special(28)
cpu.IF.instruction[13] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[14] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[15] = 32'b000000_00000_00000_00000_00000_100000;	//NOP

//special_3:
cpu.IF.instruction[16] = 32'b000000_00000_00010_10000_00000_100000;	//add r16, r0, r2
cpu.IF.instruction[17] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[18] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[19] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[20] = 32'b000000_00000_00101_01000_00000_100000;	//add r8, r0, r5
cpu.IF.instruction[21] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[22] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[23] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[24] = 32'b000010_00000_00000_00000_00011_101100;	//j print_ans(236)
cpu.IF.instruction[25] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[26] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[27] = 32'b000000_00000_00000_00000_00000_100000;	//NOP

//non_special:
cpu.IF.instruction[28] = 32'b000000_01000_00000_01001_00000_100000;	//add r9, r8, r0
cpu.IF.instruction[29] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[30] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[31] = 32'b000000_00000_00000_00000_00000_100000;	//NOP

//rem_1:
cpu.IF.instruction[32] = 32'b000000_01001_00010_01001_00000_100010;	//sub r9, r9, 2
cpu.IF.instruction[33] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[34] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[35] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[36] = 32'b000100_01001_00000_00000_00000_010111;	//beq r9, r0, even(23)
cpu.IF.instruction[37] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[38] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[39] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[40] = 32'b000100_01001_00001_00000_00000_000111;	//beq r9, r1, odd(7)
cpu.IF.instruction[41] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[42] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[43] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[44] = 32'b000010_00000_00000_00000_00000_100000;	// j rem_1(32)
cpu.IF.instruction[45] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[46] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[47] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
// odd
cpu.IF.instruction[48] = 32'b000000_01000_00010_01001_00000_100000;	//add r9, r8, r2
cpu.IF.instruction[49] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[50] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[51] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[52] = 32'b000000_01000_00010_01000_00000_100010;	//sub r8, r8, r2
cpu.IF.instruction[53] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[54] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[55] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[56] = 32'b000010_00000_00000_00000_00001_000100;	//j find_root(68)
cpu.IF.instruction[57] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[58] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[59] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
// even
cpu.IF.instruction[60] = 32'b000000_01000_00001_01001_00000_100000;	//add r9, r8, r1**
cpu.IF.instruction[61] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[62] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[63] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[64] = 32'b000000_01000_00001_01000_00000_100010;	//sub r8, r8, r1
cpu.IF.instruction[65] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[66] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[67] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
// find_root
cpu.IF.instruction[68] = 32'b000000_00000_01000_01101_00000_100000;	//add r13, r0, r8
cpu.IF.instruction[69] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[70] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[71] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[72] = 32'b000000_00000_00000_01010_00000_100000;
cpu.IF.instruction[73] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[74] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[75] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[76] = 32'b000000_00000_00001_01011_00000_100000;
cpu.IF.instruction[77] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[78] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[79] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[80] = 32'b001001_01011_01011_0000000000001111;   	//sll  _$t3, _$t3, _30    ;
cpu.IF.instruction[81] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[82] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[83] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[84] = 32'b000000_01101_01011_11000_00000_101010;
cpu.IF.instruction[85] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[86] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[87] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[88] = 32'b000100_11000_00000_00000_00000_001011;
cpu.IF.instruction[89] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[90] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[91] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[92] = 32'b001010_01011_01011_0000000000000010;   	//srl $_t3, $_t3, 2_;
cpu.IF.instruction[93] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[94] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[95] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[96] = 32'b000010_00000_00000_00000_00001_010100;
cpu.IF.instruction[97] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[98] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[99] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[100] = 32'b000100_01011_00000_00000_00000_101011;
cpu.IF.instruction[101] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[102] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[103] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[104] = 32'b000000_01010_01011_01100_00000_100000;
cpu.IF.instruction[105] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[106] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[107] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[108] = 32'b000000_01101_01100_11000_00000_101010;
cpu.IF.instruction[109] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[110] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[111] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[112] = 32'b000100_11000_00000_00000_00000_001011;
cpu.IF.instruction[113] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[114] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[115] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[116] = 32'b001010_01010_01010_0000000000000001;	 //srl $_t2, $_t2, 1_;
cpu.IF.instruction[117] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[118] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[119] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[120] = 32'b000010_00000_00000_00000_00010_001000;
cpu.IF.instruction[121] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[122] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[123] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[124] = 32'b000000_01101_01100_01101_00000_100010;
cpu.IF.instruction[125] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[126] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[127] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[128] = 32'b001010_01010_01010_0000000000000001;	 //srl $_t2, $_t2, 1_;
cpu.IF.instruction[129] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[130] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[131] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[132] = 32'b000000_01010_01011_01010_00000_100000;
cpu.IF.instruction[133] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[134] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[135] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[136] = 32'b001010_01011_01011_0000000000000010;  	//srl $_t3, $_t3, 2_;
cpu.IF.instruction[137] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[138] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[139] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[140] = 32'b000010_00000_00000_00000_00001_100100;
cpu.IF.instruction[141] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[142] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[143] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[144] = 32'b000000_00000_00011_01011_00000_100000;
cpu.IF.instruction[145] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[146] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[147] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[148] = 32'b000000_01010_01011_11000_00000_101010;
cpu.IF.instruction[149] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[150] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[151] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[152] = 32'b000100_11000_00001_00000_00000_111011;
cpu.IF.instruction[153] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[154] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[155] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[156] = 32'b000000_01000_00000_01100_00000_100000;
cpu.IF.instruction[157] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[158] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[159] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[160] = 32'b000100_01100_01011_00000_00000_011111;
cpu.IF.instruction[161] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[162] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[163] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[164] = 32'b000000_01100_01011_11001_00000_101010;
cpu.IF.instruction[165] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[166] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[167] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[168] = 32'b000100_11001_00000_00000_00000_000111;
cpu.IF.instruction[169] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[170] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[171] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[172] = 32'b000100_11001_00001_00000_00000_001011;
cpu.IF.instruction[173] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[174] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[175] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[176] = 32'b000000_01100_01011_01100_00000_100010;
cpu.IF.instruction[177] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[178] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[179] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[180] = 32'b000010_00000_00000_00000_00010_100000;
cpu.IF.instruction[181] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[182] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[183] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[184] = 32'b000000_01011_00010_01011_00000_100000;
cpu.IF.instruction[185] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[186] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[187] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[188] = 32'b000010_00000_00000_00000_00010_010100;
cpu.IF.instruction[189] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[190] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[191] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[192] = 32'b000100_10011_00001_00000_00000_001011;
cpu.IF.instruction[193] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[194] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[195] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[196] = 32'b000000_01000_00010_01000_00000_100010;
cpu.IF.instruction[197] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[198] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[199] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[200] = 32'b000010_00000_00000_00000_00001_000100;
cpu.IF.instruction[201] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[202] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[203] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[204] = 32'b000000_01000_00010_01000_00000_100000;
cpu.IF.instruction[205] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[206] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[207] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[208] = 32'b000010_00000_00000_00000_00001_000100;
cpu.IF.instruction[209] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[210] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[211] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[212] = 32'b000100_10011_00000_00000_00000_000111;
cpu.IF.instruction[213] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[214] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[215] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[216] = 32'b000100_10011_00001_00000_00000_010011;
cpu.IF.instruction[217] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[218] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[219] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[220] = 32'b000000_00000_01000_10000_00000_100000;
cpu.IF.instruction[221] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[222] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[223] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[224] = 32'b000000_00000_01001_01000_00000_100000;
cpu.IF.instruction[225] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[226] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[227] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[228] = 32'b000000_10011_00001_10011_00000_100000;
cpu.IF.instruction[229] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[230] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[231] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[232] = 32'b000010_00000_00000_00000_00001_000100;
cpu.IF.instruction[233] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[234] = 32'b000000_00000_00000_00000_00000_100000;
cpu.IF.instruction[235] = 32'b000000_00000_00000_00000_00000_100000;
// ## print_ans
cpu.IF.instruction[236] = 32'b101011_00000_01000_0000000000000001;	//sw r0, r8, 1
cpu.IF.instruction[237] = 32'b101011_00000_10000_0000000000000010;	//sw r0, r16, 2
cpu.IF.instruction[238] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[239] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
cpu.IF.instruction[240] = 32'b000000_00000_00000_00000_00000_100000;	//NOP
		
		
	for (i=241; i<300; i=i+1)  cpu.IF.instruction[ i] = 32'b000000_00000_00000_00000_00000_100000;	//NOP(add $0, $0, $0)
	cpu.IF.PC = 0;
end

//clock cycle time is 20ns, inverse Clk value per 10ns
initial Clk = 1'b1;
always #(`CYCLE_TIME/2) Clk = ~Clk;

//Rst signal
initial begin
	cycles = 32'b0;
	Rst = 1'b1;
	#12 Rst = 1'b0;
end

CPU cpu(
	.clk(Clk),
	.rst(Rst)
);

//display all Register value and Data memory content
always @(posedge Clk) begin
	cycles <= cycles + 1;
	if (cycles == `INSTRUCTION_NUMBERS) $finish; // Finish when excute the 24-th instruction (End label).
	$display("PC: %d cycles: %d", cpu.FD_PC>>2 , cycles);
	$display("  R00-R07: %08x %08x %08x %08x %08x %08x %08x %08x", cpu.ID.REG[0], cpu.ID.REG[1], cpu.ID.REG[2], cpu.ID.REG[3],cpu.ID.REG[4], cpu.ID.REG[5], cpu.ID.REG[6], cpu.ID.REG[7]);
	$display("  R08-R15: %08x %08x %08x %08x %08x %08x %08x %08x", cpu.ID.REG[8], cpu.ID.REG[9], cpu.ID.REG[10], cpu.ID.REG[11],cpu.ID.REG[12], cpu.ID.REG[13], cpu.ID.REG[14], cpu.ID.REG[15]);
	$display("  R16-R23: %08x %08x %08x %08x %08x %08x %08x %08x", cpu.ID.REG[16], cpu.ID.REG[17], cpu.ID.REG[18], cpu.ID.REG[19],cpu.ID.REG[20], cpu.ID.REG[21], cpu.ID.REG[22], cpu.ID.REG[23]);
	$display("  R24-R31: %08x %08x %08x %08x %08x %08x %08x %08x", cpu.ID.REG[24], cpu.ID.REG[25], cpu.ID.REG[26], cpu.ID.REG[27],cpu.ID.REG[28], cpu.ID.REG[29], cpu.ID.REG[30], cpu.ID.REG[31]);
	$display("  0x00   : %08x %08x %08x %08x %08x %08x %08x %08x", cpu.MEM.DM[0],cpu.MEM.DM[1],cpu.MEM.DM[2],cpu.MEM.DM[3],cpu.MEM.DM[4],cpu.MEM.DM[5],cpu.MEM.DM[6],cpu.MEM.DM[7]);
	$display("  0x08   : %08x %08x %08x %08x %08x %08x %08x %08x", cpu.MEM.DM[8],cpu.MEM.DM[9],cpu.MEM.DM[10],cpu.MEM.DM[11],cpu.MEM.DM[12],cpu.MEM.DM[13],cpu.MEM.DM[14],cpu.MEM.DM[15]);
end

//generate wave file, it can use gtkwave to display
initial begin
	$dumpfile("cpu_hw.vcd");
	$dumpvars;
end
endmodule

